//module primitive_device(
//  input clk_i,
//  input rst_i
//);

//  wire [4:0]  A1;
//  wire [4:0]  A2;
//  wire [4:0]  A3;
  
//  wire        WE3;

//  wire [31:0] RD1;
//  wire [31:0] RD2;

//  RF rf(
//    .A1( A1 ),
//    .A2( A2 ),
    

//endmodule
