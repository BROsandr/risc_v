module csr(

);
endmodule
