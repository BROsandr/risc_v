// fpga4student.com: FPGA projects, Verilog projects, VHDL projects
// FPGA tutorial: seven-segment LED display controller on Basys  3 FPGA
module Seven_segment_LED_Display_Controller(
    input clock_100Mhz, // 100 Mhz clock source on Basys 3 FPGA
    input reset, // reset
    input logic [15:0] displayed_number_i,
    
    output reg [3:0] AN, // anode signals of the 7-segment LED display
    output reg [6:0] SEG// cathode patterns of the 7-segment LED display
    );
    
//    function [15:0] to_BCD( input [13:0] bin );
   
//      integer i;
//      logic [15:0] bcd;
//      bcd=0;		 	
//      for (i=0;i<14;i=i+1) begin					//Iterate once for each bit in input number
//        if (bcd[3:0] >= 5) bcd[3:0] = bcd[3:0] + 3;		//If any BCD digit is >= 5, add three
//        if (bcd[7:4] >= 5) bcd[7:4] = bcd[7:4] + 3;
//        if (bcd[11:8] >= 5) bcd[11:8] = bcd[11:8] + 3;
//        if (bcd[15:12] >= 5) bcd[15:12] = bcd[15:12] + 3;
//        bcd = {bcd[14:0],bin[13-i]};				//Shift one bit, and shift in proper bit from input 
//      end
      
//      return bcd;
//    endfunction
    
//    assign displayed_number_i = to_BCD(32);
    
    wire rst = reset;
    
    reg [3:0]  LED_BCD;
    reg [19:0] refresh_counter; // 20-bit for creating 10.5ms refresh period or 380Hz refresh rate
             // the first 2 MSB bits for creating 4 LED-activating signals with 2.6ms digit period
    wire [1:0] LED_activating_counter; 
                 // count     0    ->  1  ->  2  ->  3
              // activates    LED1    LED2   LED3   LED4
             // and repeat        
             
    always_ff @(posedge clock_100Mhz or posedge rst)
    begin 
        if( rst==1 )
            refresh_counter <= 0;
        else
            refresh_counter <= refresh_counter + 1;
    end 
    assign LED_activating_counter = refresh_counter[19:18];
    // anode activating signals for 4 LEDs, digit period of 2.6ms
    // decoder to generate anode signals 
    always_comb
    begin
        case(LED_activating_counter)
        2'b00: begin
            AN = 4'b0111; 
            // activate LED1 and Deactivate LED2, LED3, LED4
            LED_BCD = displayed_number_i[15:12];
            // the first digit of the 16-bit number
              end
        2'b01: begin
            AN = 4'b1011; 
            // activate LED2 and Deactivate LED1, LED3, LED4
            LED_BCD = displayed_number_i[11:8];
            // the second digit of the 16-bit number
              end
        2'b10: begin
            AN = 4'b1101; 
            // activate LED3 and Deactivate LED2, LED1, LED4
            LED_BCD = displayed_number_i[7:4];
            // the third digit of the 16-bit number
                end
        2'b11: begin
            AN = 4'b1110; 
            // activate LED4 and Deactivate LED2, LED3, LED1
            LED_BCD = displayed_number_i[3:0];
            // the fourth digit of the 16-bit number    
               end
        endcase
    end
    // Cathode patterns of the 7-segment LED display 
    always_comb
    begin
        case(LED_BCD)
        4'b0000: SEG = 7'b0000001; // "0"     
        4'b0001: SEG = 7'b1001111; // "1" 
        4'b0010: SEG = 7'b0010010; // "2" 
        4'b0011: SEG = 7'b0000110; // "3" 
        4'b0100: SEG = 7'b1001100; // "4" 
        4'b0101: SEG = 7'b0100100; // "5" 
        4'b0110: SEG = 7'b0100000; // "6" 
        4'b0111: SEG = 7'b0001111; // "7" 
        4'b1000: SEG = 7'b0000000; // "8"     
        4'b1001: SEG = 7'b0000100; // "9" 
        default: SEG = 7'b0000001; // "0"
        endcase
    end
 endmodule